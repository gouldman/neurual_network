`timescale 1ns/1ps

module fake_conv_control_tb;

  // ----------------------------
  // Parameters
  // ----------------------------
  parameter WIDTH = 8;
  parameter kernel_size = 5;
  parameter pic_size = 28;
  parameter SIGN = 1;
  parameter FP_POSITIONS = 4;
  parameter channel = 3;
  parameter kernel_number = 4;

  // ----------------------------
  // Interface signals
  // ----------------------------
  logic clk;
  logic rst_n;
  logic [WIDTH-1:0] pic;
  logic pic_valid;
  logic conv_start;
  logic need_pic;
  logic conv_finish;
  logic conv_result_valid;
  logic [WIDTH-1:0] conv_result;
  logic [$clog2(pic_size*pic_size)-1:0] conv_result_addr;

  // ----------------------------
  // Clock Generation
  // ----------------------------
  initial begin
    clk = 0;
    forever #5 clk = ~clk; // 100MHz clock
  end

  // ----------------------------
  // DUT instantiation
  // ----------------------------
  fake_conv_control #(
    .WIDTH(WIDTH),
    .kernel_size(kernel_size),
    .pic_size(pic_size),
    .SIGN(SIGN),
    .FP_POSITIONS(FP_POSITIONS),
    .channel(channel),
    .kernel_number(kernel_number)
  ) dut (
    .clk(clk),
    .rst_n(rst_n),
    .pic(pic),
    .pic_valid(pic_valid),
    .conv_start(conv_start),
    .need_pic(need_pic),
    .conv_finish(conv_finish),
    .conv_result_valid(conv_result_valid),
    .conv_result(conv_result),
    .conv_result_addr(conv_result_addr)
  );

  // ----------------------------
  // Reset Task
  // ----------------------------
  task automatic reset_dut();
    begin
      rst_n = 0;
      pic = '0;
      pic_valid = 0;
      conv_start = 0;
      @(posedge clk);
      @(posedge clk);
      rst_n = 1;
      @(posedge clk);
    end
  endtask

  // ----------------------------
  // Stimulus Task
  // ----------------------------
  // ----------------------------
  // Test Sequence
  // ----------------------------
  initial begin
    reset_dut(); 
    conv_start = 1;
    #10;
    conv_start = 0;
    #100;
    pic_valid = 1;
    #100000;
        #100000;
            #100000;
                    #100000;
    $finish;
  end

endmodule

